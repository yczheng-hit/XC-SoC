module AHBlite_Decoder #(parameter Port0_en = 1,
                         parameter Port1_en = 1,
                         parameter Port2_en = 1,
                         parameter Port3_en = 1,
                         parameter Port4_en = 1)
                        (input [31:0] HADDR,
                         output wire P0_HSEL,
                         output wire P1_HSEL,
                         output wire P2_HSEL,
                         output wire P3_HSEL,
                         output wire P4_HSEL);
    
    //RAMCODE-----------------------------------
    
    //0x00000000-0x0000ffff
    /*Insert RAMCODE decoder code there*/
    assign P0_HSEL = (HADDR[31:16] == 16'h0000) ? Port0_en : 1'b0;
    /***********************************/
    
    //RAMDATA-----------------------------
    //0X20000000-0X2000FFFF
    /*Insert RAMDATA decoder code there*/
    assign P1_HSEL = (HADDR[31:16] == 16'h2000) ? Port1_en : 1'b0;
    /***********************************/
    
    //PERIPHRAL-----------------------------
    //0X40010000-0X4001FFFF
    /*Insert RAMDATA decoder code there*/
    assign P2_HSEL = (HADDR[31:16] == 16'h4001) ? Port2_en : 1'b0;
    /***********************************/
    
    //0X40000010 UART RX DATA
    //0X40000014 UART TX STATE
    //0X40000018 UART TX DATA
    /*Insert UART decoder code there*/
    assign P3_HSEL = (HADDR[31:4] == 28'h4000001) ? Port3_en : 1'b0;
    /***********************************/
    
    assign P4_HSEL = (HADDR[31:4] == 28'h4000002) ? Port4_en : 1'b0;
    
endmodule
